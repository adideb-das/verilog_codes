module and_gate(
    //Input and Output Parameters
    input wire a,
    input wire b,
    output wire y
);

//and gate function
assign y = a & b;

endmodule
