module or_gate(
    //Input and Output Parameters
    input wire a,
    input wire b,
    output wire y
);
//or gate function
assign y = a | b;

endmodule